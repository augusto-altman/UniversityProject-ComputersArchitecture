`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:16:38 05/27/2014 
// Design Name: 
// Module Name:    ControlHazzardHandler 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ControlHazzardHandler(
    input isJump,
    output reg stall_exe,
    output reg stall_id
    );

	
	
endmodule
